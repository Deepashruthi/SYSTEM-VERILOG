// DYNAMIC ARRAY ORDERING
module dynamic_array2;
  int array[] = '{1,6,4,3,5};
  initial begin
    $display("size = %0d",array.size());
    array.reverse();
    $display(array);
    array.sort();
    $display(array);
    array.rsort();
    $display(array);
    array.shuffle();
    $display(array);
  end
endmodule
