//Interface
interface inter;
  logic clk;
  logic rst;
  logic u_d;
  logic [3:0] count;
endinterface
