//Interface
interface inter();
  logic clk;
  logic rst;
  logic d;
  logic q;
endinterface
