//Interface 
interface inter();
  logic clk;
  logic wr;
  logic [7:0] data_i;
  logic [7:0] data_o;
  logic [3:0] addr;
endinterface
